module CONTROLUNIT( 

AR_LOAD, AR_INC, 
PC_BUS, PC_LOAD, PC_INC,
DR_BUS_H, DR_BUS_L, DR_LOAD,
TR_BUS, TR_LOAD,
IR_LOAD,
R_BUS, R_LOAD,
AC_BUS, AC_LOAD,
ALUS7, ALUS6, ALUS5, ALUS4, ALUS3, ALUS2, ALUS1,
Z_LOAD,

MEMBUS, BUSMEM, WE,

IR, CLK, CLEAR, INC, Z);

input IR, CLK, CLEAR, INC, Z;

output AR_LOAD, AR_INC, 
PC_BUS, PC_LOAD, PC_INC,
DR_BUS_H, DR_BUS_L, DR_LOAD,
TR_BUS, TR_LOAD,
IR_LOAD,
R_BUS, R_LOAD,
AC_BUS, AC_LOAD,
ALUS7, ALUS6, ALUS5, ALUS4, ALUS3, ALUS2, ALUS1,
Z_LOAD,
MEMBUS, BUSMEM, WE;

CONTROL_COMB CU_COMB( 

AR_LOAD, AR_INC, 
PC_BUS, PC_LOAD, PC_INC,
DR_BUS_H, DR_BUS_L, DR_LOAD,
TR_BUS, TR_LOAD,
IR_LOAD,
R_BUS, R_LOAD,
AC_BUS, AC_LOAD,
ALUS7, ALUS6, ALUS5, ALUS4, ALUS3, ALUS2, ALUS1,
Z_LOAD,

MEMBUS, BUSMEM, WE,
IR, CLK, CLEAR, INC, Z);

endmodule 
