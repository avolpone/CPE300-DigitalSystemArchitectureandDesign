module AC(AC_OUT, BUS, AC_BUS, Z_LOAD, AC_LOAD, CLK);

	output reg [7:0] AC_OUT; 

	input [7:0] BUS; 

	input CLK, AC_LOAD, Z_LOAD, AC_BUS;
	
	reg [7:0] AC_temp, Z;
	
	wire [7:0] ALU_OUT, ZCHECKED;
	
ALU ALUMOD(ALU_OUT, ALUS7, ALUS6, ALUS5, ALUS4, ALUS3, ALUS2, ALUS1, BUS, AC_temp);	

Z_CHECK ZCHECK(ZCHECKED, Z_LOAD, ALU_OUT);

always
	Z = ZCHECKED;

always @(posedge CLK)
begin
	if(AC_LOAD)
		AC_temp <= ALU_OUT;
	else if(!AC_LOAD)
		AC_temp <= AC_temp;
end
	
always
begin
	if(AC_BUS)
		AC_OUT <= AC_temp;
	else if(!AC_BUS)
		AC_OUT = 8'bz;
end
	
endmodule 