module CENTRAL_PROCESSOR(AC_TOCPU, PC_TOCPU, CLK, START, FULL_RESET);

input CLK, START, FULL_RESET;

output [7:0] AC_TOCPU;
output [15:0] PC_TOCPU;

wire
INCREMENT,
CLOCK_ENABLED,
COUNT_RESET, 
SOFT_RESET,

AR_LOAD, AR_INC, 
PC_BUS, PC_LOAD, PC_INC, PC_RESET,
DR_BUS_H, DR_BUS_L, DR_LOAD,
TR_BUS, TR_LOAD,
IR_LOAD,
R_BUS, R_LOAD,
AC_BUS, AC_LOAD,
ALUS7, ALUS6, ALUS5, ALUS4, ALUS3, ALUS2, ALUS1,
Z_LOAD,

MEMBUS, BUSMEM, WE,

IR, CLK, CLEAR, INC, Z, Z_TOCU;

wire [7:0] IR_TOCU;

and (CLOCK_ENABLED, CLK, START);
or(INCREMENT, START, FULL_RESET);

CONTROL_STEP CONTROLSTEP( T0, T1, T2, T3, T4, T5, T6, T7, INCREMENT,
INOP, ILDAC, ISTAC, IMVAC, IMOVR, IJUMP, IJMPZ, IJPNZ, IADD, ISUB, IINAC, ICLAC, IAND, IOR, IXOR, INOT, IR_TOCU, 
SOFT_RESET, FULL_RESET, CLOCK_ENABLED);

CONTROL_COMB CU( SOFT_RESET,

AR_LOAD, AR_INC, 
PC_BUS, PC_LOAD, PC_INC, PC_RESET,
DR_BUS_H, DR_BUS_L, DR_LOAD,
TR_BUS, TR_LOAD,
IR_LOAD,
R_BUS, R_LOAD,
AC_BUS, AC_LOAD,
ALUS7, ALUS6, ALUS5, ALUS4, ALUS3, ALUS2, ALUS1,

MEMBUS, BUSMEM, WE,

T0, T1, T2, T3, T4, T5, T6, T7,
INOP, ILDAC, ISTAC, IMVAC, IMOVR, IJUMP, IJMPZ, IJPNZ, IADD, ISUB, IINAC, ICLAC, IAND, IOR, IXOR, INOT, FULL_RESET, Z_TOCU);

DATAPATH DP( PC_TOCPU, AC_TOCPU, IR_TOCU, Z_TOCU,
AR_LOAD, AR_INC, 
PC_BUS, PC_LOAD, PC_INC, PC_RESET,
DR_BUS_H, DR_BUS_L, DR_LOAD,
TR_BUS, TR_LOAD,
IR_LOAD,
R_BUS, R_LOAD,
AC_BUS, AC_LOAD,
ALUS7, ALUS6, ALUS5, ALUS4, ALUS3, ALUS2, ALUS1,

MEMBUS, BUSMEM, WE, CLOCK_ENABLED);

assign IR_TOCPU = IR_TOCU;

/*
BCD_8bit BCD(AC_TOCPU, HUNDREDS, TENS, ONES);
sevenseg oneseg(ONES, AC_ONES);
sevenseg tenseg(TENS, AC_TENS);
sevenseg hunseg(HUNDREDS, AC_HUNDREDS);
*/
endmodule 
